module pc_update (
    input clk,
    input p_cnd,
    input [3:0] D_icode,
    input [63:0] D_valC,
    input [63:0] D_valP,

    output reg F_PC
);
    

endmodule