module and_64b(
  input signed [63:0]a,
  input signed [63:0]b,
  output signed [63:0]out
);

genvar i;
generate
    for(i=0;i<64;i=i+1)begin
    and g1 (out[i],a[i],b[i]);
    end
endgenerate

endmodule

